module webp

pub enum AlphaFilter {
	@none
	fast
	best
}
