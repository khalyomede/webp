module webp

pub struct Resize {
	width int = 0
	height int = 0
}
