module webp

pub enum Metadata {
	all
	@none
	exif
	icc
	xmp
}
