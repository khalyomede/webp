module webp

pub enum Preset {
	@none
	_default
	photo
	picture
	drawing
	icon
	text
}
