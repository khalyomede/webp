module webp

pub struct Crop {
	x_position int [required]
	y_position int [required]
	width int [required]
	height int [required]
}
