module webp

pub enum Hint {
	@none
	photo
	picture
	graph
}
